//Modulo que permite convertir se?ales logicas de distintos niveles de tensi?n
//De momento esta versi?n no tiene entradas bididreccionales, pero se puede intentar(TODO)



module level_shifter (
    input  VIN, //se?al de entrada 
    input  VCC_LOW, //fuente de alimentaci?n de nivel bajo
    input  VCC_HIGH, //fuente de alimentaci?n de nivel alto
    output real VOUT //se?al de salida 

    );

 

endmodule
